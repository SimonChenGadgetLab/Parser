
Signal a : std_logic_vector (0 to 3);
signal b : std_logic_vector(0 to 2);
signal C : std_logic; 


if (a = b) then a <= c; elsif (a < c) then a <= b else	
if (a = b) then
		a <= '0' & '1' & b(1 downto 0);
	        b <= (others => '0');  
	        --b <= (others => '1');
		if (c = 4)
		c <=B"1111"; 

			--abc
